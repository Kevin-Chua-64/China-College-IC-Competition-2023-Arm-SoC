
module BUFG (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
